`timescale 1ns/1ns
module MSDFF(input D, clk, rst, output Q, Qb);