`timescale 1ns/1ns

module TB_s10000001detector;
    reg clk, rst, J;
    wire Y;
        s10000001detectorQ DUT (.clk(clk), .rst(rst), .J(J), .Y(Y));

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
        rst = 1;
        J = 0;
        #20;
        rst = 0;
        #20;

        J = 0; #10;
        J = 1; #10;
        J = 0; #10;
        J = 0; #10;
        J = 1; #10;
        J = 0; #10;
        J = 1; #10;

        J = 1; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 1; #10;

        J = 1; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 1; #10;
        J = 0; #10;

        J = 0; #10;
        J = 1; #10;
        J = 1; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;

        J = 1; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 0; #10;
        J = 1; #10;

        #50;
        $stop;
    end

endmodule

