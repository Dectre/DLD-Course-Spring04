`timescale 1ns/1ns
module TB_6();
logic [1:0] A, B;
wire g;
function_g cutG(A, B, g);
initial begin
for (int i = 0; i < 4; i++) begin
for (int j = 0; j < 4; j++) begin
A = i[1:0];
B = j[1:0];
#271;
end
end
end
endmodule;

