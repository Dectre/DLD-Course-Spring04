`timescale 1ns/1ns
module myOAI_switch(input a, b, c, output w);
supply1 vdd; supply0 gnd;
wire i,j;
pmos #(5, 6, 7) T1(i, vdd, a), T2(w, i, b), T3(w, vdd, c);
nmos #(3, 4, 5) T4(j, gnd, a), T5(j, gnd, b), T6(w, j, c);
endmodule
